Preemp Test Netlist
.INCLUDE constants.cir
.INCLUDE popamp.cir
.INCLUDE hp.cir
.INCLUDE lp.cir
.INCLUDE gain.cir
.INCLUDE preemp.cir
Vin	0	1	AC	1
Xpe	1	2	preemp
.AC DEC 40 100 10k
.PRINT VDB(2)
.options list
.options post
.END
