.SUBCKT	pgain in out
* K=27.67dB
Rf	n	out	24.2k
Ri	in	n	1k
X1	0	n	out	popamp
.ENDS pgain
