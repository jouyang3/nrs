Summing Op-Amp Test
.INCLUDE popamp.cir
.INCLUDE sum.cir

V1	0	1	1
V2	0	2	1
Xs	1	2	out	sum

.TRAN	100NS	1us
.PRINT	v(out)
.OPTION POST
.END
