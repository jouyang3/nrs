.SUBCKT joint in out
X1	in	out	out	popamp
.ENDS joint