Test

.SUBCKT popamp 	4 	n 	2
Ri	4	n	2MEG
Ei	1	0	4	n	1
R	1	3	1
C	3	0	0.03183
Eo	6	0	3	0	200K
Ro	6	2	75
.ENDS popamp

.SUBCKT php in out
C1	in	1	1
R1	1	out	0.707
C2	1	p	1
R2	p	0	1.414
X1	p	out	out	popamp
.ENDS php

.SUBCKT plp in out
R1	in	1	1
R2	1	p	1
C1	1	out	1.414
C2	p	0	0.707
X1	p	out	out
.ENDS plp

.SUBCKT	pgain in out
Rf	n	out	15.8
Ri	in	n	1
X1	0	n	out	popamp
.ENDS pgain

.SUBCKT preemp in out
Xhp	in	1	php
Xlp	1	2	plp
Xg	2	out	pgain
.ENDS preemp

Vin	0	1	AC	1
Xpe	1	2	preemp
R1	2	0	1K


.AC DEC 40 100 10K
.PRINT VDB(2), VP(2)
.OPTIONS POST
.END
