.PARAM Pi=3.1415926535897932384626433832795028841971693993751058
