.SUBCKT preemp in out
.PARAM khf='2*500*Pi'
.PARAM klf='w0^2/khf'
Xhp	in	1	hp	kf=khf	c=2n
Xlp	1	2	lp	kf=klf	r=120k
Xg	2	out	gain	a='10^(29/20)'
.ENDS preemp
