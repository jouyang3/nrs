Preemphasis Gain
.SUBCKT	pgain in out
Rf	n	out	15.8
Ri	in	n	1
X1	0	n	out	popamp
.ENDS pgain