.SUBCKT php in out
C1	in	1	2n
R1	1	out	112523
C2	1	p	2n
R2	p	0	225045
X1	p	out	out	popamp
.ENDS php
