.SUBCKT sum 