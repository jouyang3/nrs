Preemphasis Low Pass
.SUBCKT plp in out
R1	in	1	1
R2	1	p	1
C1	1	out	1.414
C2	p	0	0.707
X1	p	out	out
.ENDS plp